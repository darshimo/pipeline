`timescale 1ns / 100ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 2016/09/08 14:33:18
// Design Name:
// Module Name: char_rom
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module char_rom(
    rst,
    addr,
    dout
    );
    input rst;
    input [10:0] addr;
    output [7:0] dout;

    reg [7:0] ch_rom [0:2047];

    assign dout = ch_rom[addr];

    always @(posedge rst) begin
        if(rst) begin
//0
            ch_rom[0] <= 8'h00;
            ch_rom[1] <= 8'h00;
            ch_rom[2] <= 8'h00;
            ch_rom[3] <= 8'h00;
            ch_rom[4] <= 8'h00;
            ch_rom[5] <= 8'h00;
            ch_rom[6] <= 8'h00;
            ch_rom[7] <= 8'h00;
            ch_rom[8] <= 8'h00;
//1
            ch_rom[9] <= 8'h00;
            ch_rom[10] <= 8'h00;
            ch_rom[11] <= 8'h00;
            ch_rom[12] <= 8'h00;
            ch_rom[13] <= 8'h00;
            ch_rom[14] <= 8'h00;
            ch_rom[15] <= 8'h00;
            ch_rom[16] <= 8'h00;
//2
            ch_rom[17] <= 8'h00;
            ch_rom[18] <= 8'h00;
            ch_rom[19] <= 8'h00;
            ch_rom[20] <= 8'h00;
            ch_rom[21] <= 8'h00;
            ch_rom[22] <= 8'h00;
            ch_rom[23] <= 8'h00;
            ch_rom[24] <= 8'h00;
//3
            ch_rom[25] <= 8'h00;
            ch_rom[26] <= 8'h00;
            ch_rom[27] <= 8'h00;
            ch_rom[28] <= 8'h00;
            ch_rom[29] <= 8'h00;
            ch_rom[30] <= 8'h00;
            ch_rom[31] <= 8'h00;
            ch_rom[32] <= 8'h00;
//4
            ch_rom[33] <= 8'h00;
            ch_rom[34] <= 8'h00;
            ch_rom[35] <= 8'h00;
            ch_rom[36] <= 8'h00;
            ch_rom[37] <= 8'h00;
            ch_rom[38] <= 8'h00;
            ch_rom[39] <= 8'h00;
            ch_rom[40] <= 8'h00;
//5
            ch_rom[41] <= 8'h00;
            ch_rom[42] <= 8'h00;
            ch_rom[43] <= 8'h00;
            ch_rom[44] <= 8'h00;
            ch_rom[45] <= 8'h00;
            ch_rom[46] <= 8'h00;
            ch_rom[47] <= 8'h00;
            ch_rom[48] <= 8'h00;
//6
            ch_rom[49] <= 8'h00;
            ch_rom[50] <= 8'h00;
            ch_rom[51] <= 8'h00;
            ch_rom[52] <= 8'h00;
            ch_rom[53] <= 8'h00;
            ch_rom[54] <= 8'h00;
            ch_rom[55] <= 8'h00;
            ch_rom[56] <= 8'h00;
//7
            ch_rom[57] <= 8'h00;
            ch_rom[58] <= 8'h00;
            ch_rom[59] <= 8'h00;
            ch_rom[60] <= 8'h00;
            ch_rom[61] <= 8'h00;
            ch_rom[62] <= 8'h00;
            ch_rom[63] <= 8'h00;
            ch_rom[64] <= 8'h00;
//8
            ch_rom[65] <= 8'h00;
            ch_rom[66] <= 8'h00;
            ch_rom[67] <= 8'h00;
            ch_rom[68] <= 8'h00;
            ch_rom[69] <= 8'h00;
            ch_rom[70] <= 8'h00;
            ch_rom[71] <= 8'h00;
            ch_rom[72] <= 8'h00;
//9
            ch_rom[73] <= 8'h00;
            ch_rom[74] <= 8'h00;
            ch_rom[75] <= 8'h00;
            ch_rom[76] <= 8'h00;
            ch_rom[77] <= 8'h00;
            ch_rom[78] <= 8'h00;
            ch_rom[79] <= 8'h00;
            ch_rom[80] <= 8'h00;
//A
            ch_rom[81] <= 8'h00;
            ch_rom[82] <= 8'h00;
            ch_rom[83] <= 8'h00;
            ch_rom[84] <= 8'h00;
            ch_rom[85] <= 8'h00;
            ch_rom[86] <= 8'h00;
            ch_rom[87] <= 8'h00;
            ch_rom[88] <= 8'h00;
//B
            ch_rom[89] <= 8'h00;
            ch_rom[90] <= 8'h00;
            ch_rom[91] <= 8'h00;
            ch_rom[92] <= 8'h00;
            ch_rom[93] <= 8'h00;
            ch_rom[94] <= 8'h00;
            ch_rom[95] <= 8'h00;
            ch_rom[96] <= 8'h00;
//C
            ch_rom[97] <= 8'h00;
            ch_rom[98] <= 8'h00;
            ch_rom[99] <= 8'h00;
            ch_rom[100] <= 8'h00;
            ch_rom[101] <= 8'h00;
            ch_rom[102] <= 8'h00;
            ch_rom[103] <= 8'h00;
            ch_rom[104] <= 8'h00;
//D
            ch_rom[105] <= 8'h00;
            ch_rom[106] <= 8'h00;
            ch_rom[107] <= 8'h00;
            ch_rom[108] <= 8'h00;
            ch_rom[109] <= 8'h00;
            ch_rom[110] <= 8'h00;
            ch_rom[111] <= 8'h00;
            ch_rom[112] <= 8'h00;
//E
            ch_rom[113] <= 8'h00;
            ch_rom[114] <= 8'h00;
            ch_rom[115] <= 8'h00;
            ch_rom[116] <= 8'h00;
            ch_rom[117] <= 8'h00;
            ch_rom[118] <= 8'h00;
            ch_rom[119] <= 8'h00;
            ch_rom[120] <= 8'h00;
//F
            ch_rom[121] <= 8'h00;
            ch_rom[122] <= 8'h00;
            ch_rom[123] <= 8'h00;
            ch_rom[124] <= 8'h00;
            ch_rom[125] <= 8'h00;
            ch_rom[126] <= 8'h00;
            ch_rom[127] <= 8'h00;
            ch_rom[128] <= 8'h00;
//10
            ch_rom[129] <= 8'h00;
            ch_rom[130] <= 8'h00;
            ch_rom[131] <= 8'h00;
            ch_rom[132] <= 8'h00;
            ch_rom[133] <= 8'h00;
            ch_rom[134] <= 8'h00;
            ch_rom[135] <= 8'h00;
            ch_rom[136] <= 8'h00;
//11
            ch_rom[137] <= 8'h00;
            ch_rom[138] <= 8'h00;
            ch_rom[139] <= 8'h00;
            ch_rom[140] <= 8'h00;
            ch_rom[141] <= 8'h00;
            ch_rom[142] <= 8'h00;
            ch_rom[143] <= 8'h00;
            ch_rom[144] <= 8'h00;
//12
            ch_rom[145] <= 8'h00;
            ch_rom[146] <= 8'h00;
            ch_rom[147] <= 8'h00;
            ch_rom[148] <= 8'h00;
            ch_rom[149] <= 8'h00;
            ch_rom[150] <= 8'h00;
            ch_rom[151] <= 8'h00;
            ch_rom[152] <= 8'h00;
//13
            ch_rom[153] <= 8'h00;
            ch_rom[154] <= 8'h00;
            ch_rom[155] <= 8'h00;
            ch_rom[156] <= 8'h00;
            ch_rom[157] <= 8'h00;
            ch_rom[158] <= 8'h00;
            ch_rom[159] <= 8'h00;
            ch_rom[160] <= 8'h00;
//14
            ch_rom[161] <= 8'h00;
            ch_rom[162] <= 8'h00;
            ch_rom[163] <= 8'h00;
            ch_rom[164] <= 8'h00;
            ch_rom[165] <= 8'h00;
            ch_rom[166] <= 8'h00;
            ch_rom[167] <= 8'h00;
            ch_rom[168] <= 8'h00;
//15
            ch_rom[169] <= 8'h00;
            ch_rom[170] <= 8'h00;
            ch_rom[171] <= 8'h00;
            ch_rom[172] <= 8'h00;
            ch_rom[173] <= 8'h00;
            ch_rom[174] <= 8'h00;
            ch_rom[175] <= 8'h00;
            ch_rom[176] <= 8'h00;
//16
            ch_rom[177] <= 8'h00;
            ch_rom[178] <= 8'h00;
            ch_rom[179] <= 8'h00;
            ch_rom[180] <= 8'h00;
            ch_rom[181] <= 8'h00;
            ch_rom[182] <= 8'h00;
            ch_rom[183] <= 8'h00;
            ch_rom[184] <= 8'h00;
//17
            ch_rom[185] <= 8'h00;
            ch_rom[186] <= 8'h00;
            ch_rom[187] <= 8'h00;
            ch_rom[188] <= 8'h00;
            ch_rom[189] <= 8'h00;
            ch_rom[190] <= 8'h00;
            ch_rom[191] <= 8'h00;
            ch_rom[192] <= 8'h00;
//18
            ch_rom[193] <= 8'h00;
            ch_rom[194] <= 8'h00;
            ch_rom[195] <= 8'h00;
            ch_rom[196] <= 8'h00;
            ch_rom[197] <= 8'h00;
            ch_rom[198] <= 8'h00;
            ch_rom[199] <= 8'h00;
            ch_rom[200] <= 8'h00;
//19
            ch_rom[201] <= 8'h00;
            ch_rom[202] <= 8'h00;
            ch_rom[203] <= 8'h00;
            ch_rom[204] <= 8'h00;
            ch_rom[205] <= 8'h00;
            ch_rom[206] <= 8'h00;
            ch_rom[207] <= 8'h00;
            ch_rom[208] <= 8'h00;
//1A
            ch_rom[209] <= 8'h00;
            ch_rom[210] <= 8'h00;
            ch_rom[211] <= 8'h00;
            ch_rom[212] <= 8'h00;
            ch_rom[213] <= 8'h00;
            ch_rom[214] <= 8'h00;
            ch_rom[215] <= 8'h00;
            ch_rom[216] <= 8'h00;
//1B
            ch_rom[217] <= 8'h00;
            ch_rom[218] <= 8'h00;
            ch_rom[219] <= 8'h00;
            ch_rom[220] <= 8'h00;
            ch_rom[221] <= 8'h00;
            ch_rom[222] <= 8'h00;
            ch_rom[223] <= 8'h00;
            ch_rom[224] <= 8'h00;
//1C
            ch_rom[225] <= 8'h00;
            ch_rom[226] <= 8'h00;
            ch_rom[227] <= 8'h00;
            ch_rom[228] <= 8'h00;
            ch_rom[229] <= 8'h00;
            ch_rom[230] <= 8'h00;
            ch_rom[231] <= 8'h00;
            ch_rom[232] <= 8'h00;
//1D
            ch_rom[233] <= 8'h00;
            ch_rom[234] <= 8'h00;
            ch_rom[235] <= 8'h00;
            ch_rom[236] <= 8'h00;
            ch_rom[237] <= 8'h00;
            ch_rom[238] <= 8'h00;
            ch_rom[239] <= 8'h00;
            ch_rom[240] <= 8'h00;
//1E
            ch_rom[241] <= 8'h00;
            ch_rom[242] <= 8'h00;
            ch_rom[243] <= 8'h00;
            ch_rom[244] <= 8'h00;
            ch_rom[245] <= 8'h00;
            ch_rom[246] <= 8'h00;
            ch_rom[247] <= 8'h00;
            ch_rom[248] <= 8'h00;
//1F
            ch_rom[249] <= 8'h00;
            ch_rom[250] <= 8'h00;
            ch_rom[251] <= 8'h00;
            ch_rom[252] <= 8'h00;
            ch_rom[253] <= 8'h00;
            ch_rom[254] <= 8'h00;
            ch_rom[255] <= 8'h00;
            ch_rom[256] <= 8'h00;
//20
            ch_rom[257] <= 8'h00;
            ch_rom[258] <= 8'h00;
            ch_rom[259] <= 8'h00;
            ch_rom[260] <= 8'h00;
            ch_rom[261] <= 8'h00;
            ch_rom[262] <= 8'h00;
            ch_rom[263] <= 8'h00;
            ch_rom[264] <= 8'h00;
//21 !
            ch_rom[265] <= 8'h00;
            ch_rom[266] <= 8'h00;
            ch_rom[267] <= 8'h5f;
            ch_rom[268] <= 8'h00;
            ch_rom[269] <= 8'h00;
            ch_rom[270] <= 8'h00;
            ch_rom[271] <= 8'h00;
            ch_rom[272] <= 8'h00;
//22 "
            ch_rom[273] <= 8'h00;
            ch_rom[274] <= 8'h03;
            ch_rom[275] <= 8'h00;
            ch_rom[276] <= 8'h03;
            ch_rom[277] <= 8'h00;
            ch_rom[278] <= 8'h00;
            ch_rom[279] <= 8'h00;
            ch_rom[280] <= 8'h64;
//23 #
            ch_rom[281] <= 8'h3c;
            ch_rom[282] <= 8'h26;
            ch_rom[283] <= 8'h64;
            ch_rom[284] <= 8'h3c;
            ch_rom[285] <= 8'h26;
            ch_rom[286] <= 8'h24;
            ch_rom[287] <= 8'h00;
            ch_rom[288] <= 8'h26;
//24 $
            ch_rom[289] <= 8'h49;
            ch_rom[290] <= 8'h49;
            ch_rom[291] <= 8'h7f;
            ch_rom[292] <= 8'h49;
            ch_rom[293] <= 8'h49;
            ch_rom[294] <= 8'h32;
            ch_rom[295] <= 8'h00;
            ch_rom[296] <= 8'h42;
//25 %
            ch_rom[297] <= 8'h25;
            ch_rom[298] <= 8'h12;
            ch_rom[299] <= 8'h08;
            ch_rom[300] <= 8'h24;
            ch_rom[301] <= 8'h52;
            ch_rom[302] <= 8'h21;
            ch_rom[303] <= 8'h00;
            ch_rom[304] <= 8'h20;
//26 &
            ch_rom[305] <= 8'h50;
            ch_rom[306] <= 8'h4e;
            ch_rom[307] <= 8'h55;
            ch_rom[308] <= 8'h22;
            ch_rom[309] <= 8'h58;
            ch_rom[310] <= 8'h28;
            ch_rom[311] <= 8'h00;
            ch_rom[312] <= 8'h00;
//27 '
            ch_rom[313] <= 8'h00;
            ch_rom[314] <= 8'h00;
            ch_rom[315] <= 8'h03;
            ch_rom[316] <= 8'h00;
            ch_rom[317] <= 8'h00;
            ch_rom[318] <= 8'h00;
            ch_rom[319] <= 8'h00;
            ch_rom[320] <= 8'h00;
//28 (
            ch_rom[321] <= 8'h00;
            ch_rom[322] <= 8'h1c;
            ch_rom[323] <= 8'h22;
            ch_rom[324] <= 8'h41;
            ch_rom[325] <= 8'h00;
            ch_rom[326] <= 8'h00;
            ch_rom[327] <= 8'h00;
            ch_rom[328] <= 8'h00;
//29 )
            ch_rom[329] <= 8'h00;
            ch_rom[330] <= 8'h00;
            ch_rom[331] <= 8'h41;
            ch_rom[332] <= 8'h22;
            ch_rom[333] <= 8'h1c;
            ch_rom[334] <= 8'h00;
            ch_rom[335] <= 8'h00;
            ch_rom[336] <= 8'h00;
//2A *
            ch_rom[337] <= 8'h15;
            ch_rom[338] <= 8'h15;
            ch_rom[339] <= 8'h0e;
            ch_rom[340] <= 8'h0e;
            ch_rom[341] <= 8'h15;
            ch_rom[342] <= 8'h15;
            ch_rom[343] <= 8'h00;
            ch_rom[344] <= 8'h00;
//2B +
            ch_rom[345] <= 8'h08;
            ch_rom[346] <= 8'h08;
            ch_rom[347] <= 8'h3e;
            ch_rom[348] <= 8'h08;
            ch_rom[349] <= 8'h08;
            ch_rom[350] <= 8'h00;
            ch_rom[351] <= 8'h00;
            ch_rom[352] <= 8'h00;
//2C ,
            ch_rom[353] <= 8'h00;
            ch_rom[354] <= 8'h00;
            ch_rom[355] <= 8'h50;
            ch_rom[356] <= 8'h30;
            ch_rom[357] <= 8'h00;
            ch_rom[358] <= 8'h00;
            ch_rom[359] <= 8'h00;
            ch_rom[360] <= 8'h00;
//2D -
            ch_rom[361] <= 8'h08;
            ch_rom[362] <= 8'h08;
            ch_rom[363] <= 8'h08;
            ch_rom[364] <= 8'h08;
            ch_rom[365] <= 8'h08;
            ch_rom[366] <= 8'h00;
            ch_rom[367] <= 8'h00;
            ch_rom[368] <= 8'h00;
//2E .
            ch_rom[369] <= 8'h00;
            ch_rom[370] <= 8'h00;
            ch_rom[371] <= 8'h40;
            ch_rom[372] <= 8'h00;
            ch_rom[373] <= 8'h00;
            ch_rom[374] <= 8'h00;
            ch_rom[375] <= 8'h00;
            ch_rom[376] <= 8'h40;
//2F /
            ch_rom[377] <= 8'h20;
            ch_rom[378] <= 8'h10;
            ch_rom[379] <= 8'h08;
            ch_rom[380] <= 8'h04;
            ch_rom[381] <= 8'h02;
            ch_rom[382] <= 8'h01;
            ch_rom[383] <= 8'h00;
            ch_rom[384] <= 8'h00;
//30 0
            ch_rom[385] <= 8'h3e;
            ch_rom[386] <= 8'h41;
            ch_rom[387] <= 8'h41;
            ch_rom[388] <= 8'h41;
            ch_rom[389] <= 8'h3e;
            ch_rom[390] <= 8'h00;
            ch_rom[391] <= 8'h00;
            ch_rom[392] <= 8'h00;
//31 1
            ch_rom[393] <= 8'h00;
            ch_rom[394] <= 8'h41;
            ch_rom[395] <= 8'h7f;
            ch_rom[396] <= 8'h40;
            ch_rom[397] <= 8'h00;
            ch_rom[398] <= 8'h00;
            ch_rom[399] <= 8'h00;
            ch_rom[400] <= 8'h00;
//32 2
            ch_rom[401] <= 8'h42;
            ch_rom[402] <= 8'h61;
            ch_rom[403] <= 8'h51;
            ch_rom[404] <= 8'h49;
            ch_rom[405] <= 8'h6e;
            ch_rom[406] <= 8'h00;
            ch_rom[407] <= 8'h00;
            ch_rom[408] <= 8'h00;
//33 3
            ch_rom[409] <= 8'h22;
            ch_rom[410] <= 8'h41;
            ch_rom[411] <= 8'h49;
            ch_rom[412] <= 8'h49;
            ch_rom[413] <= 8'h36;
            ch_rom[414] <= 8'h00;
            ch_rom[415] <= 8'h00;
            ch_rom[416] <= 8'h00;
//34 4
            ch_rom[417] <= 8'h18;
            ch_rom[418] <= 8'h14;
            ch_rom[419] <= 8'h12;
            ch_rom[420] <= 8'h7f;
            ch_rom[421] <= 8'h10;
            ch_rom[422] <= 8'h00;
            ch_rom[423] <= 8'h00;
            ch_rom[424] <= 8'h00;
//35 5
            ch_rom[425] <= 8'h27;
            ch_rom[426] <= 8'h49;
            ch_rom[427] <= 8'h49;
            ch_rom[428] <= 8'h49;
            ch_rom[429] <= 8'h71;
            ch_rom[430] <= 8'h00;
            ch_rom[431] <= 8'h00;
            ch_rom[432] <= 8'h00;
//36 6
            ch_rom[433] <= 8'h3c;
            ch_rom[434] <= 8'h4a;
            ch_rom[435] <= 8'h49;
            ch_rom[436] <= 8'h48;
            ch_rom[437] <= 8'h70;
            ch_rom[438] <= 8'h00;
            ch_rom[439] <= 8'h00;
            ch_rom[440] <= 8'h00;
//37 7
            ch_rom[441] <= 8'h43;
            ch_rom[442] <= 8'h21;
            ch_rom[443] <= 8'h11;
            ch_rom[444] <= 8'h0d;
            ch_rom[445] <= 8'h03;
            ch_rom[446] <= 8'h00;
            ch_rom[447] <= 8'h00;
            ch_rom[448] <= 8'h00;
//38 8
            ch_rom[449] <= 8'h36;
            ch_rom[450] <= 8'h49;
            ch_rom[451] <= 8'h49;
            ch_rom[452] <= 8'h49;
            ch_rom[453] <= 8'h36;
            ch_rom[454] <= 8'h00;
            ch_rom[455] <= 8'h00;
            ch_rom[456] <= 8'h00;
//39 9
            ch_rom[457] <= 8'h06;
            ch_rom[458] <= 8'h09;
            ch_rom[459] <= 8'h49;
            ch_rom[460] <= 8'h29;
            ch_rom[461] <= 8'h1e;
            ch_rom[462] <= 8'h00;
            ch_rom[463] <= 8'h00;
            ch_rom[464] <= 8'h00;
//3a
            ch_rom[465] <= 8'h00;
            ch_rom[466] <= 8'h00;
            ch_rom[467] <= 8'h12;
            ch_rom[468] <= 8'h00;
            ch_rom[469] <= 8'h00;
            ch_rom[470] <= 8'h00;
            ch_rom[471] <= 8'h00;
            ch_rom[472] <= 8'h00;
//3b
            ch_rom[473] <= 8'h00;
            ch_rom[474] <= 8'h00;
            ch_rom[475] <= 8'h52;
            ch_rom[476] <= 8'h30;
            ch_rom[477] <= 8'h00;
            ch_rom[478] <= 8'h00;
            ch_rom[479] <= 8'h00;
            ch_rom[480] <= 8'h00;
//3c
            ch_rom[481] <= 8'h00;
            ch_rom[482] <= 8'h08;
            ch_rom[483] <= 8'h14;
            ch_rom[484] <= 8'h14;
            ch_rom[485] <= 8'h22;
            ch_rom[486] <= 8'h00;
            ch_rom[487] <= 8'h00;
            ch_rom[488] <= 8'h00;
//3d
            ch_rom[489] <= 8'h14;
            ch_rom[490] <= 8'h14;
            ch_rom[491] <= 8'h14;
            ch_rom[492] <= 8'h14;
            ch_rom[493] <= 8'h14;
            ch_rom[494] <= 8'h14;
            ch_rom[495] <= 8'h00;
            ch_rom[496] <= 8'h00;
//3e
            ch_rom[497] <= 8'h00;
            ch_rom[498] <= 8'h22;
            ch_rom[499] <= 8'h14;
            ch_rom[500] <= 8'h14;
            ch_rom[501] <= 8'h08;
            ch_rom[502] <= 8'h00;
            ch_rom[503] <= 8'h00;
            ch_rom[504] <= 8'h00;
//3f
            ch_rom[505] <= 8'h02;
            ch_rom[506] <= 8'h01;
            ch_rom[507] <= 8'h59;
            ch_rom[508] <= 8'h05;
            ch_rom[509] <= 8'h02;
            ch_rom[510] <= 8'h00;
            ch_rom[511] <= 8'h00;
            ch_rom[512] <= 8'h3e;
//40
            ch_rom[513] <= 8'h41;
            ch_rom[514] <= 8'h5d;
            ch_rom[515] <= 8'h55;
            ch_rom[516] <= 8'h4d;
            ch_rom[517] <= 8'h51;
            ch_rom[518] <= 8'h2e;
            ch_rom[519] <= 8'h00;
            ch_rom[520] <= 8'h40;
//41 A
            ch_rom[521] <= 8'h7c;
            ch_rom[522] <= 8'h4a;
            ch_rom[523] <= 8'h09;
            ch_rom[524] <= 8'h4a;
            ch_rom[525] <= 8'h7c;
            ch_rom[526] <= 8'h40;
            ch_rom[527] <= 8'h00;
            ch_rom[528] <= 8'h41;
//42 B
            ch_rom[529] <= 8'h7f;
            ch_rom[530] <= 8'h49;
            ch_rom[531] <= 8'h49;
            ch_rom[532] <= 8'h49;
            ch_rom[533] <= 8'h49;
            ch_rom[534] <= 8'h36;
            ch_rom[535] <= 8'h00;
            ch_rom[536] <= 8'h1c;
//43 C
            ch_rom[537] <= 8'h22;
            ch_rom[538] <= 8'h41;
            ch_rom[539] <= 8'h41;
            ch_rom[540] <= 8'h41;
            ch_rom[541] <= 8'h41;
            ch_rom[542] <= 8'h22;
            ch_rom[543] <= 8'h00;
            ch_rom[544] <= 8'h41;
//44 D
            ch_rom[545] <= 8'h7f;
            ch_rom[546] <= 8'h41;
            ch_rom[547] <= 8'h41;
            ch_rom[548] <= 8'h41;
            ch_rom[549] <= 8'h22;
            ch_rom[550] <= 8'h1c;
            ch_rom[551] <= 8'h00;
            ch_rom[552] <= 8'h41;
//45 E
            ch_rom[553] <= 8'h7f;
            ch_rom[554] <= 8'h49;
            ch_rom[555] <= 8'h49;
            ch_rom[556] <= 8'h5d;
            ch_rom[557] <= 8'h41;
            ch_rom[558] <= 8'h63;
            ch_rom[559] <= 8'h00;
            ch_rom[560] <= 8'h41;
//46 F
            ch_rom[561] <= 8'h7f;
            ch_rom[562] <= 8'h49;
            ch_rom[563] <= 8'h09;
            ch_rom[564] <= 8'h1d;
            ch_rom[565] <= 8'h01;
            ch_rom[566] <= 8'h03;
            ch_rom[567] <= 8'h00;
            ch_rom[568] <= 8'h1c;
//47 G
            ch_rom[569] <= 8'h22;
            ch_rom[570] <= 8'h41;
            ch_rom[571] <= 8'h49;
            ch_rom[572] <= 8'h49;
            ch_rom[573] <= 8'h3a;
            ch_rom[574] <= 8'h08;
            ch_rom[575] <= 8'h00;
            ch_rom[576] <= 8'h41;
//48 H
            ch_rom[577] <= 8'h7f;
            ch_rom[578] <= 8'h08;
            ch_rom[579] <= 8'h08;
            ch_rom[580] <= 8'h08;
            ch_rom[581] <= 8'h7f;
            ch_rom[582] <= 8'h41;
            ch_rom[583] <= 8'h00;
            ch_rom[584] <= 8'h00;
//49 I
            ch_rom[585] <= 8'h41;
            ch_rom[586] <= 8'h41;
            ch_rom[587] <= 8'h7F;
            ch_rom[588] <= 8'h41;
            ch_rom[589] <= 8'h41;
            ch_rom[590] <= 8'h00;
            ch_rom[591] <= 8'h00;
            ch_rom[592] <= 8'h30;
//4A J
            ch_rom[593] <= 8'h40;
            ch_rom[594] <= 8'h41;
            ch_rom[595] <= 8'h41;
            ch_rom[596] <= 8'h3F;
            ch_rom[597] <= 8'h01;
            ch_rom[598] <= 8'h01;
            ch_rom[599] <= 8'h00;
            ch_rom[600] <= 8'h41;
//4B K
            ch_rom[601] <= 8'h7f;
            ch_rom[602] <= 8'h08;
            ch_rom[603] <= 8'h0c;
            ch_rom[604] <= 8'h12;
            ch_rom[605] <= 8'h61;
            ch_rom[606] <= 8'h41;
            ch_rom[607] <= 8'h00;
            ch_rom[608] <= 8'h41;
//4C L
            ch_rom[609] <= 8'h7f;
            ch_rom[610] <= 8'h41;
            ch_rom[611] <= 8'h40;
            ch_rom[612] <= 8'h40;
            ch_rom[613] <= 8'h40;
            ch_rom[614] <= 8'h60;
            ch_rom[615] <= 8'h00;
            ch_rom[616] <= 8'h41;
//4D M
            ch_rom[617] <= 8'h7f;
            ch_rom[618] <= 8'h42;
            ch_rom[619] <= 8'h0c;
            ch_rom[620] <= 8'h42;
            ch_rom[621] <= 8'h7f;
            ch_rom[622] <= 8'h41;
            ch_rom[623] <= 8'h00;
            ch_rom[624] <= 8'h41;
//4E N
            ch_rom[625] <= 8'h7f;
            ch_rom[626] <= 8'h42;
            ch_rom[627] <= 8'h0c;
            ch_rom[628] <= 8'h11;
            ch_rom[629] <= 8'h7f;
            ch_rom[630] <= 8'h01;
            ch_rom[631] <= 8'h00;
            ch_rom[632] <= 8'h1c;
//4F O
            ch_rom[633] <= 8'h22;
            ch_rom[634] <= 8'h41;
            ch_rom[635] <= 8'h41;
            ch_rom[636] <= 8'h41;
            ch_rom[637] <= 8'h22;
            ch_rom[638] <= 8'h1c;
            ch_rom[639] <= 8'h00;
            ch_rom[640] <= 8'h41;
//50 P
            ch_rom[641] <= 8'h7f;
            ch_rom[642] <= 8'h49;
            ch_rom[643] <= 8'h09;
            ch_rom[644] <= 8'h09;
            ch_rom[645] <= 8'h09;
            ch_rom[646] <= 8'h06;
            ch_rom[647] <= 8'h00;
            ch_rom[648] <= 8'h0c;
//51 Q
            ch_rom[649] <= 8'h12;
            ch_rom[650] <= 8'h21;
            ch_rom[651] <= 8'h21;
            ch_rom[652] <= 8'h61;
            ch_rom[653] <= 8'h52;
            ch_rom[654] <= 8'h4c;
            ch_rom[655] <= 8'h00;
            ch_rom[656] <= 8'h41;
//52 R
            ch_rom[657] <= 8'h7f;
            ch_rom[658] <= 8'h09;
            ch_rom[659] <= 8'h09;
            ch_rom[660] <= 8'h19;
            ch_rom[661] <= 8'h69;
            ch_rom[662] <= 8'h46;
            ch_rom[663] <= 8'h00;
            ch_rom[664] <= 8'h66;
//53 S
            ch_rom[665] <= 8'h49;
            ch_rom[666] <= 8'h49;
            ch_rom[667] <= 8'h49;
            ch_rom[668] <= 8'h49;
            ch_rom[669] <= 8'h49;
            ch_rom[670] <= 8'h33;
            ch_rom[671] <= 8'h00;
            ch_rom[672] <= 8'h03;
//54 T
            ch_rom[673] <= 8'h01;
            ch_rom[674] <= 8'h41;
            ch_rom[675] <= 8'h7f;
            ch_rom[676] <= 8'h41;
            ch_rom[677] <= 8'h01;
            ch_rom[678] <= 8'h03;
            ch_rom[679] <= 8'h00;
            ch_rom[680] <= 8'h01;
//55 U
            ch_rom[681] <= 8'h3f;
            ch_rom[682] <= 8'h41;
            ch_rom[683] <= 8'h40;
            ch_rom[684] <= 8'h41;
            ch_rom[685] <= 8'h3f;
            ch_rom[686] <= 8'h01;
            ch_rom[687] <= 8'h00;
            ch_rom[688] <= 8'h01;
//56 V
            ch_rom[689] <= 8'h0f;
            ch_rom[690] <= 8'h31;
            ch_rom[691] <= 8'h40;
            ch_rom[692] <= 8'h31;
            ch_rom[693] <= 8'h0f;
            ch_rom[694] <= 8'h01;
            ch_rom[695] <= 8'h00;
            ch_rom[696] <= 8'h01;
//57 W
            ch_rom[697] <= 8'h1f;
            ch_rom[698] <= 8'h61;
            ch_rom[699] <= 8'h14;
            ch_rom[700] <= 8'h61;
            ch_rom[701] <= 8'h1f;
            ch_rom[702] <= 8'h01;
            ch_rom[703] <= 8'h00;
            ch_rom[704] <= 8'h41;
//58 X
            ch_rom[705] <= 8'h41;
            ch_rom[706] <= 8'h36;
            ch_rom[707] <= 8'h08;
            ch_rom[708] <= 8'h36;
            ch_rom[709] <= 8'h41;
            ch_rom[710] <= 8'h41;
            ch_rom[711] <= 8'h00;
            ch_rom[712] <= 8'h01;
//59 Y
            ch_rom[713] <= 8'h03;
            ch_rom[714] <= 8'h44;
            ch_rom[715] <= 8'h78;
            ch_rom[716] <= 8'h44;
            ch_rom[717] <= 8'h03;
            ch_rom[718] <= 8'h01;
            ch_rom[719] <= 8'h00;
            ch_rom[720] <= 8'h43;
//5A Z
            ch_rom[721] <= 8'h61;
            ch_rom[722] <= 8'h51;
            ch_rom[723] <= 8'h49;
            ch_rom[724] <= 8'h45;
            ch_rom[725] <= 8'h43;
            ch_rom[726] <= 8'h61;
            ch_rom[727] <= 8'h00;
            ch_rom[728] <= 8'h00;
//5B
            ch_rom[729] <= 8'h00;
            ch_rom[730] <= 8'h7f;
            ch_rom[731] <= 8'h41;
            ch_rom[732] <= 8'h41;
            ch_rom[733] <= 8'h00;
            ch_rom[734] <= 8'h00;
            ch_rom[735] <= 8'h00;
            ch_rom[736] <= 8'h01;
//5C
            ch_rom[737] <= 8'h02;
            ch_rom[738] <= 8'h04;
            ch_rom[739] <= 8'h08;
            ch_rom[740] <= 8'h10;
            ch_rom[741] <= 8'h20;
            ch_rom[742] <= 8'h40;
            ch_rom[743] <= 8'h00;
            ch_rom[744] <= 8'h00;
//5D
            ch_rom[745] <= 8'h00;
            ch_rom[746] <= 8'h41;
            ch_rom[747] <= 8'h41;
            ch_rom[748] <= 8'h7f;
            ch_rom[749] <= 8'h00;
            ch_rom[750] <= 8'h00;
            ch_rom[751] <= 8'h00;
            ch_rom[752] <= 8'h00;
//5E
            ch_rom[753] <= 8'h04;
            ch_rom[754] <= 8'h02;
            ch_rom[755] <= 8'h01;
            ch_rom[756] <= 8'h01;
            ch_rom[757] <= 8'h02;
            ch_rom[758] <= 8'h04;
            ch_rom[759] <= 8'h00;
            ch_rom[760] <= 8'h00;
//5F
            ch_rom[761] <= 8'h40;
            ch_rom[762] <= 8'h40;
            ch_rom[763] <= 8'h40;
            ch_rom[764] <= 8'h40;
            ch_rom[765] <= 8'h40;
            ch_rom[766] <= 8'h40;
            ch_rom[767] <= 8'h00;
            ch_rom[768] <= 8'h00;
//60
            ch_rom[769] <= 8'h01;
            ch_rom[770] <= 8'h02;
            ch_rom[771] <= 8'h00;
            ch_rom[772] <= 8'h00;
            ch_rom[773] <= 8'h00;
            ch_rom[774] <= 8'h00;
            ch_rom[775] <= 8'h00;
            ch_rom[776] <= 8'h00;
//61 a
            ch_rom[777] <= 8'h34;
            ch_rom[778] <= 8'h4a;
            ch_rom[779] <= 8'h4a;
            ch_rom[780] <= 8'h4a;
            ch_rom[781] <= 8'h3c;
            ch_rom[782] <= 8'h40;
            ch_rom[783] <= 8'h00;
            ch_rom[784] <= 8'h00;
//62 b
            ch_rom[785] <= 8'h41;
            ch_rom[786] <= 8'h3f;
            ch_rom[787] <= 8'h48;
            ch_rom[788] <= 8'h48;
            ch_rom[789] <= 8'h48;
            ch_rom[790] <= 8'h30;
            ch_rom[791] <= 8'h00;
            ch_rom[792] <= 8'h00;
//63 c
            ch_rom[793] <= 8'h3c;
            ch_rom[794] <= 8'h42;
            ch_rom[795] <= 8'h42;
            ch_rom[796] <= 8'h42;
            ch_rom[797] <= 8'h24;
            ch_rom[798] <= 8'h00;
            ch_rom[799] <= 8'h00;
            ch_rom[800] <= 8'h00;
//64 d
            ch_rom[801] <= 8'h30;
            ch_rom[802] <= 8'h48;
            ch_rom[803] <= 8'h48;
            ch_rom[804] <= 8'h49;
            ch_rom[805] <= 8'h3f;
            ch_rom[806] <= 8'h40;
            ch_rom[807] <= 8'h00;
            ch_rom[808] <= 8'h00;
//65 e
            ch_rom[809] <= 8'h3c;
            ch_rom[810] <= 8'h4a;
            ch_rom[811] <= 8'h4a;
            ch_rom[812] <= 8'h4a;
            ch_rom[813] <= 8'h2c;
            ch_rom[814] <= 8'h00;
            ch_rom[815] <= 8'h00;
            ch_rom[816] <= 8'h00;
//66 f
            ch_rom[817] <= 8'h00;
            ch_rom[818] <= 8'h48;
            ch_rom[819] <= 8'h7e;
            ch_rom[820] <= 8'h49;
            ch_rom[821] <= 8'h09;
            ch_rom[822] <= 8'h00;
            ch_rom[823] <= 8'h00;
            ch_rom[824] <= 8'h00;
//67 g
            ch_rom[825] <= 8'h26;
            ch_rom[826] <= 8'h49;
            ch_rom[827] <= 8'h49;
            ch_rom[828] <= 8'h49;
            ch_rom[829] <= 8'h3f;
            ch_rom[830] <= 8'h01;
            ch_rom[831] <= 8'h00;
            ch_rom[832] <= 8'h41;
//68 h
            ch_rom[833] <= 8'h7f;
            ch_rom[834] <= 8'h48;
            ch_rom[835] <= 8'h04;
            ch_rom[836] <= 8'h44;
            ch_rom[837] <= 8'h78;
            ch_rom[838] <= 8'h40;
            ch_rom[839] <= 8'h00;
            ch_rom[840] <= 8'h00;
//69 i
            ch_rom[841] <= 8'h00;
            ch_rom[842] <= 8'h44;
            ch_rom[843] <= 8'h7d;
            ch_rom[844] <= 8'h40;
            ch_rom[845] <= 8'h00;
            ch_rom[846] <= 8'h00;
            ch_rom[847] <= 8'h00;
            ch_rom[848] <= 8'h00;
//6a j
            ch_rom[849] <= 8'h00;
            ch_rom[850] <= 8'h40;
            ch_rom[851] <= 8'h44;
            ch_rom[852] <= 8'h3d;
            ch_rom[853] <= 8'h00;
            ch_rom[854] <= 8'h00;
            ch_rom[855] <= 8'h00;
            ch_rom[856] <= 8'h41;
//6b k
            ch_rom[857] <= 8'h7f;
            ch_rom[858] <= 8'h10;
            ch_rom[859] <= 8'h18;
            ch_rom[860] <= 8'h24;
            ch_rom[861] <= 8'h42;
            ch_rom[862] <= 8'h42;
            ch_rom[863] <= 8'h00;
            ch_rom[864] <= 8'h00;
//6c l
            ch_rom[865] <= 8'h40;
            ch_rom[866] <= 8'h41;
            ch_rom[867] <= 8'h7f;
            ch_rom[868] <= 8'h40;
            ch_rom[869] <= 8'h40;
            ch_rom[870] <= 8'h00;
            ch_rom[871] <= 8'h00;
            ch_rom[872] <= 8'h42;
//6d m
            ch_rom[873] <= 8'h7e;
            ch_rom[874] <= 8'h02;
            ch_rom[875] <= 8'h7c;
            ch_rom[876] <= 8'h02;
            ch_rom[877] <= 8'h7e;
            ch_rom[878] <= 8'h40;
            ch_rom[879] <= 8'h00;
            ch_rom[880] <= 8'h42;
//6e n
            ch_rom[881] <= 8'h7e;
            ch_rom[882] <= 8'h44;
            ch_rom[883] <= 8'h02;
            ch_rom[884] <= 8'h42;
            ch_rom[885] <= 8'h7c;
            ch_rom[886] <= 8'h40;
            ch_rom[887] <= 8'h00;
            ch_rom[888] <= 8'h00;
//6f o
            ch_rom[889] <= 8'h3c;
            ch_rom[890] <= 8'h42;
            ch_rom[891] <= 8'h42;
            ch_rom[892] <= 8'h42;
            ch_rom[893] <= 8'h3c;
            ch_rom[894] <= 8'h00;
            ch_rom[895] <= 8'h00;
            ch_rom[896] <= 8'h00;
//70 p
            ch_rom[897] <= 8'h41;
            ch_rom[898] <= 8'h7f;
            ch_rom[899] <= 8'h49;
            ch_rom[900] <= 8'h09;
            ch_rom[901] <= 8'h09;
            ch_rom[902] <= 8'h06;
            ch_rom[903] <= 8'h00;
            ch_rom[904] <= 8'h00;
//71 q
            ch_rom[905] <= 8'h06;
            ch_rom[906] <= 8'h09;
            ch_rom[907] <= 8'h09;
            ch_rom[908] <= 8'h49;
            ch_rom[909] <= 8'h7f;
            ch_rom[910] <= 8'h41;
            ch_rom[911] <= 8'h00;
            ch_rom[912] <= 8'h00;
//72 r
            ch_rom[913] <= 8'h42;
            ch_rom[914] <= 8'h7e;
            ch_rom[915] <= 8'h44;
            ch_rom[916] <= 8'h02;
            ch_rom[917] <= 8'h02;
            ch_rom[918] <= 8'h04;
            ch_rom[919] <= 8'h00;
            ch_rom[920] <= 8'h00;
//73 s
            ch_rom[921] <= 8'h64;
            ch_rom[922] <= 8'h4a;
            ch_rom[923] <= 8'h4a;
            ch_rom[924] <= 8'h4a;
            ch_rom[925] <= 8'h36;
            ch_rom[926] <= 8'h00;
            ch_rom[927] <= 8'h00;
            ch_rom[928] <= 8'h00;
//74 t
            ch_rom[929] <= 8'h04;
            ch_rom[930] <= 8'h3f;
            ch_rom[931] <= 8'h44;
            ch_rom[932] <= 8'h44;
            ch_rom[933] <= 8'h20;
            ch_rom[934] <= 8'h00;
            ch_rom[935] <= 8'h00;
            ch_rom[936] <= 8'h00;
//75 u
            ch_rom[937] <= 8'h02;
            ch_rom[938] <= 8'h3e;
            ch_rom[939] <= 8'h40;
            ch_rom[940] <= 8'h40;
            ch_rom[941] <= 8'h22;
            ch_rom[942] <= 8'h7e;
            ch_rom[943] <= 8'h40;
            ch_rom[944] <= 8'h02;
//76 v
            ch_rom[945] <= 8'h0e;
            ch_rom[946] <= 8'h32;
            ch_rom[947] <= 8'h40;
            ch_rom[948] <= 8'h32;
            ch_rom[949] <= 8'h0e;
            ch_rom[950] <= 8'h02;
            ch_rom[951] <= 8'h00;
            ch_rom[952] <= 8'h02;
//77 w
            ch_rom[953] <= 8'h1e;
            ch_rom[954] <= 8'h62;
            ch_rom[955] <= 8'h18;
            ch_rom[956] <= 8'h62;
            ch_rom[957] <= 8'h1e;
            ch_rom[958] <= 8'h02;
            ch_rom[959] <= 8'h00;
            ch_rom[960] <= 8'h42;
//78 x
            ch_rom[961] <= 8'h62;
            ch_rom[962] <= 8'h14;
            ch_rom[963] <= 8'h08;
            ch_rom[964] <= 8'h14;
            ch_rom[965] <= 8'h62;
            ch_rom[966] <= 8'h42;
            ch_rom[967] <= 8'h00;
            ch_rom[968] <= 8'h01;
//79 y
            ch_rom[969] <= 8'h43;
            ch_rom[970] <= 8'h45;
            ch_rom[971] <= 8'h38;
            ch_rom[972] <= 8'h05;
            ch_rom[973] <= 8'h03;
            ch_rom[974] <= 8'h01;
            ch_rom[975] <= 8'h00;
            ch_rom[976] <= 8'h00;
//7a z
            ch_rom[977] <= 8'h46;
            ch_rom[978] <= 8'h62;
            ch_rom[979] <= 8'h52;
            ch_rom[980] <= 8'h4a;
            ch_rom[981] <= 8'h46;
            ch_rom[982] <= 8'h62;
            ch_rom[983] <= 8'h00;
            ch_rom[984] <= 8'h00;
//7b
            ch_rom[985] <= 8'h00;
            ch_rom[986] <= 8'h08;
            ch_rom[987] <= 8'h36;
            ch_rom[988] <= 8'h41;
            ch_rom[989] <= 8'h00;
            ch_rom[990] <= 8'h00;
            ch_rom[991] <= 8'h00;
            ch_rom[992] <= 8'h00;
//7c
            ch_rom[993] <= 8'h00;
            ch_rom[994] <= 8'h00;
            ch_rom[995] <= 8'h7f;
            ch_rom[996] <= 8'h00;
            ch_rom[997] <= 8'h00;
            ch_rom[998] <= 8'h00;
            ch_rom[999] <= 8'h00;
            ch_rom[1000] <= 8'h00;
//7d
            ch_rom[1001] <= 8'h00;
            ch_rom[1002] <= 8'h00;
            ch_rom[1003] <= 8'h41;
            ch_rom[1004] <= 8'h36;
            ch_rom[1005] <= 8'h08;
            ch_rom[1006] <= 8'h00;
            ch_rom[1007] <= 8'h00;
            ch_rom[1008] <= 8'h00;
//7e
            ch_rom[1009] <= 8'h18;
            ch_rom[1010] <= 8'h08;
            ch_rom[1011] <= 8'h08;
            ch_rom[1012] <= 8'h10;
            ch_rom[1013] <= 8'h10;
            ch_rom[1014] <= 8'h18;
            ch_rom[1015] <= 8'h00;
            ch_rom[1016] <= 8'hAA;
//7f
            ch_rom[1017] <= 8'h55;
            ch_rom[1018] <= 8'hAA;
            ch_rom[1019] <= 8'h55;
            ch_rom[1020] <= 8'hAA;
            ch_rom[1021] <= 8'h55;
            ch_rom[1022] <= 8'hAA;
            ch_rom[1023] <= 8'h55;

            ch_rom[1024] <= 8'h00;
            ch_rom[1025] <= 8'h00;
            ch_rom[1026] <= 8'h00;
            ch_rom[1027] <= 8'h00;
            ch_rom[1028] <= 8'h00;
            ch_rom[1029] <= 8'h00;
            ch_rom[1030] <= 8'h00;
            ch_rom[1031] <= 8'h00;
            ch_rom[1032] <= 8'h00;
            ch_rom[1033] <= 8'h00;
            ch_rom[1034] <= 8'h00;
            ch_rom[1035] <= 8'h00;
            ch_rom[1036] <= 8'h00;
            ch_rom[1037] <= 8'h00;
            ch_rom[1038] <= 8'h00;
            ch_rom[1039] <= 8'h00;
            ch_rom[1040] <= 8'h00;
            ch_rom[1041] <= 8'h00;
            ch_rom[1042] <= 8'h00;
            ch_rom[1043] <= 8'h00;
            ch_rom[1044] <= 8'h00;
            ch_rom[1045] <= 8'h00;
            ch_rom[1046] <= 8'h00;
            ch_rom[1047] <= 8'h00;
            ch_rom[1048] <= 8'h00;
            ch_rom[1049] <= 8'h00;
            ch_rom[1050] <= 8'h00;
            ch_rom[1051] <= 8'h00;
            ch_rom[1052] <= 8'h00;
            ch_rom[1053] <= 8'h00;
            ch_rom[1054] <= 8'h00;
            ch_rom[1055] <= 8'h00;
            ch_rom[1056] <= 8'h00;
            ch_rom[1057] <= 8'h00;
            ch_rom[1058] <= 8'h00;
            ch_rom[1059] <= 8'h00;
            ch_rom[1060] <= 8'h00;
            ch_rom[1061] <= 8'h00;
            ch_rom[1062] <= 8'h00;
            ch_rom[1063] <= 8'h00;
            ch_rom[1064] <= 8'h00;
            ch_rom[1065] <= 8'h00;
            ch_rom[1066] <= 8'h00;
            ch_rom[1067] <= 8'h00;
            ch_rom[1068] <= 8'h00;
            ch_rom[1069] <= 8'h00;
            ch_rom[1070] <= 8'h00;
            ch_rom[1071] <= 8'h00;
            ch_rom[1072] <= 8'h00;
            ch_rom[1073] <= 8'h00;
            ch_rom[1074] <= 8'h00;
            ch_rom[1075] <= 8'h00;
            ch_rom[1076] <= 8'h00;
            ch_rom[1077] <= 8'h00;
            ch_rom[1078] <= 8'h00;
            ch_rom[1079] <= 8'h00;
            ch_rom[1080] <= 8'h00;
            ch_rom[1081] <= 8'h00;
            ch_rom[1082] <= 8'h00;
            ch_rom[1083] <= 8'h00;
            ch_rom[1084] <= 8'h00;
            ch_rom[1085] <= 8'h00;
            ch_rom[1086] <= 8'h00;
            ch_rom[1087] <= 8'h00;
            ch_rom[1088] <= 8'h00;
            ch_rom[1089] <= 8'h00;
            ch_rom[1090] <= 8'h00;
            ch_rom[1091] <= 8'h00;
            ch_rom[1092] <= 8'h00;
            ch_rom[1093] <= 8'h00;
            ch_rom[1094] <= 8'h00;
            ch_rom[1095] <= 8'h00;
            ch_rom[1096] <= 8'h00;
            ch_rom[1097] <= 8'h00;
            ch_rom[1098] <= 8'h00;
            ch_rom[1099] <= 8'h00;
            ch_rom[1100] <= 8'h00;
            ch_rom[1101] <= 8'h00;
            ch_rom[1102] <= 8'h00;
            ch_rom[1103] <= 8'h00;
            ch_rom[1104] <= 8'h00;
            ch_rom[1105] <= 8'h00;
            ch_rom[1106] <= 8'h00;
            ch_rom[1107] <= 8'h00;
            ch_rom[1108] <= 8'h00;
            ch_rom[1109] <= 8'h00;
            ch_rom[1110] <= 8'h00;
            ch_rom[1111] <= 8'h00;
            ch_rom[1112] <= 8'h00;
            ch_rom[1113] <= 8'h00;
            ch_rom[1114] <= 8'h00;
            ch_rom[1115] <= 8'h00;
            ch_rom[1116] <= 8'h00;
            ch_rom[1117] <= 8'h00;
            ch_rom[1118] <= 8'h00;
            ch_rom[1119] <= 8'h00;
            ch_rom[1120] <= 8'h00;
            ch_rom[1121] <= 8'h00;
            ch_rom[1122] <= 8'h00;
            ch_rom[1123] <= 8'h00;
            ch_rom[1124] <= 8'h00;
            ch_rom[1125] <= 8'h00;
            ch_rom[1126] <= 8'h00;
            ch_rom[1127] <= 8'h00;
            ch_rom[1128] <= 8'h00;
            ch_rom[1129] <= 8'h00;
            ch_rom[1130] <= 8'h00;
            ch_rom[1131] <= 8'h00;
            ch_rom[1132] <= 8'h00;
            ch_rom[1133] <= 8'h00;
            ch_rom[1134] <= 8'h00;
            ch_rom[1135] <= 8'h00;
            ch_rom[1136] <= 8'h00;
            ch_rom[1137] <= 8'h00;
            ch_rom[1138] <= 8'h00;
            ch_rom[1139] <= 8'h00;
            ch_rom[1140] <= 8'h00;
            ch_rom[1141] <= 8'h00;
            ch_rom[1142] <= 8'h00;
            ch_rom[1143] <= 8'h00;
            ch_rom[1144] <= 8'h00;
            ch_rom[1145] <= 8'h00;
            ch_rom[1146] <= 8'h00;
            ch_rom[1147] <= 8'h00;
            ch_rom[1148] <= 8'h00;
            ch_rom[1149] <= 8'h00;
            ch_rom[1150] <= 8'h00;
            ch_rom[1151] <= 8'h00;
            ch_rom[1152] <= 8'h00;
            ch_rom[1153] <= 8'h00;
            ch_rom[1154] <= 8'h00;
            ch_rom[1155] <= 8'h00;
            ch_rom[1156] <= 8'h00;
            ch_rom[1157] <= 8'h00;
            ch_rom[1158] <= 8'h00;
            ch_rom[1159] <= 8'h00;
            ch_rom[1160] <= 8'h00;
            ch_rom[1161] <= 8'h00;
            ch_rom[1162] <= 8'h00;
            ch_rom[1163] <= 8'h00;
            ch_rom[1164] <= 8'h00;
            ch_rom[1165] <= 8'h00;
            ch_rom[1166] <= 8'h00;
            ch_rom[1167] <= 8'h00;
            ch_rom[1168] <= 8'h00;
            ch_rom[1169] <= 8'h00;
            ch_rom[1170] <= 8'h00;
            ch_rom[1171] <= 8'h00;
            ch_rom[1172] <= 8'h00;
            ch_rom[1173] <= 8'h00;
            ch_rom[1174] <= 8'h00;
            ch_rom[1175] <= 8'h00;
            ch_rom[1176] <= 8'h00;
            ch_rom[1177] <= 8'h00;
            ch_rom[1178] <= 8'h00;
            ch_rom[1179] <= 8'h00;
            ch_rom[1180] <= 8'h00;
            ch_rom[1181] <= 8'h00;
            ch_rom[1182] <= 8'h00;
            ch_rom[1183] <= 8'h00;
            ch_rom[1184] <= 8'h00;
            ch_rom[1185] <= 8'h00;
            ch_rom[1186] <= 8'h00;
            ch_rom[1187] <= 8'h00;
            ch_rom[1188] <= 8'h00;
            ch_rom[1189] <= 8'h00;
            ch_rom[1190] <= 8'h00;
            ch_rom[1191] <= 8'h00;
            ch_rom[1192] <= 8'h00;
            ch_rom[1193] <= 8'h00;
            ch_rom[1194] <= 8'h00;
            ch_rom[1195] <= 8'h00;
            ch_rom[1196] <= 8'h00;
            ch_rom[1197] <= 8'h00;
            ch_rom[1198] <= 8'h00;
            ch_rom[1199] <= 8'h00;
            ch_rom[1200] <= 8'h00;
            ch_rom[1201] <= 8'h00;
            ch_rom[1202] <= 8'h00;
            ch_rom[1203] <= 8'h00;
            ch_rom[1204] <= 8'h00;
            ch_rom[1205] <= 8'h00;
            ch_rom[1206] <= 8'h00;
            ch_rom[1207] <= 8'h00;
            ch_rom[1208] <= 8'h00;
            ch_rom[1209] <= 8'h00;
            ch_rom[1210] <= 8'h00;
            ch_rom[1211] <= 8'h00;
            ch_rom[1212] <= 8'h00;
            ch_rom[1213] <= 8'h00;
            ch_rom[1214] <= 8'h00;
            ch_rom[1215] <= 8'h00;
            ch_rom[1216] <= 8'h00;
            ch_rom[1217] <= 8'h00;
            ch_rom[1218] <= 8'h00;
            ch_rom[1219] <= 8'h00;
            ch_rom[1220] <= 8'h00;
            ch_rom[1221] <= 8'h00;
            ch_rom[1222] <= 8'h00;
            ch_rom[1223] <= 8'h00;
            ch_rom[1224] <= 8'h00;
            ch_rom[1225] <= 8'h00;
            ch_rom[1226] <= 8'h00;
            ch_rom[1227] <= 8'h00;
            ch_rom[1228] <= 8'h00;
            ch_rom[1229] <= 8'h00;
            ch_rom[1230] <= 8'h00;
            ch_rom[1231] <= 8'h00;
            ch_rom[1232] <= 8'h00;
            ch_rom[1233] <= 8'h00;
            ch_rom[1234] <= 8'h00;
            ch_rom[1235] <= 8'h00;
            ch_rom[1236] <= 8'h00;
            ch_rom[1237] <= 8'h00;
            ch_rom[1238] <= 8'h00;
            ch_rom[1239] <= 8'h00;
            ch_rom[1240] <= 8'h00;
            ch_rom[1241] <= 8'h00;
            ch_rom[1242] <= 8'h00;
            ch_rom[1243] <= 8'h00;
            ch_rom[1244] <= 8'h00;
            ch_rom[1245] <= 8'h00;
            ch_rom[1246] <= 8'h00;
            ch_rom[1247] <= 8'h00;
            ch_rom[1248] <= 8'h00;
            ch_rom[1249] <= 8'h00;
            ch_rom[1250] <= 8'h00;
            ch_rom[1251] <= 8'h00;
            ch_rom[1252] <= 8'h00;
            ch_rom[1253] <= 8'h00;
            ch_rom[1254] <= 8'h00;
            ch_rom[1255] <= 8'h00;
            ch_rom[1256] <= 8'h00;
            ch_rom[1257] <= 8'h00;
            ch_rom[1258] <= 8'h00;
            ch_rom[1259] <= 8'h00;
            ch_rom[1260] <= 8'h00;
            ch_rom[1261] <= 8'h00;
            ch_rom[1262] <= 8'h00;
            ch_rom[1263] <= 8'h00;
            ch_rom[1264] <= 8'h00;
            ch_rom[1265] <= 8'h00;
            ch_rom[1266] <= 8'h00;
            ch_rom[1267] <= 8'h00;
            ch_rom[1268] <= 8'h00;
            ch_rom[1269] <= 8'h00;
            ch_rom[1270] <= 8'h00;
            ch_rom[1271] <= 8'h00;
            ch_rom[1272] <= 8'h00;
            ch_rom[1273] <= 8'h00;
            ch_rom[1274] <= 8'h00;
            ch_rom[1275] <= 8'h00;
            ch_rom[1276] <= 8'h00;
            ch_rom[1277] <= 8'h00;
            ch_rom[1278] <= 8'h00;
            ch_rom[1279] <= 8'h00;
            ch_rom[1280] <= 8'h00;
            ch_rom[1281] <= 8'h00;
            ch_rom[1282] <= 8'h00;
            ch_rom[1283] <= 8'h00;
            ch_rom[1284] <= 8'h00;
            ch_rom[1285] <= 8'h00;
            ch_rom[1286] <= 8'h00;
            ch_rom[1287] <= 8'h00;
            ch_rom[1288] <= 8'h00;
            ch_rom[1289] <= 8'h00;
            ch_rom[1290] <= 8'h00;
            ch_rom[1291] <= 8'h00;
            ch_rom[1292] <= 8'h00;
            ch_rom[1293] <= 8'h00;
            ch_rom[1294] <= 8'h00;
            ch_rom[1295] <= 8'h00;
            ch_rom[1296] <= 8'h00;
            ch_rom[1297] <= 8'h00;
            ch_rom[1298] <= 8'h00;
            ch_rom[1299] <= 8'h00;
            ch_rom[1300] <= 8'h00;
            ch_rom[1301] <= 8'h00;
            ch_rom[1302] <= 8'h00;
            ch_rom[1303] <= 8'h00;
            ch_rom[1304] <= 8'h00;
            ch_rom[1305] <= 8'h00;
            ch_rom[1306] <= 8'h00;
            ch_rom[1307] <= 8'h00;
            ch_rom[1308] <= 8'h00;
            ch_rom[1309] <= 8'h00;
            ch_rom[1310] <= 8'h00;
            ch_rom[1311] <= 8'h00;
            ch_rom[1312] <= 8'h00;
            ch_rom[1313] <= 8'h00;
            ch_rom[1314] <= 8'h00;
            ch_rom[1315] <= 8'h00;
            ch_rom[1316] <= 8'h00;
            ch_rom[1317] <= 8'h00;
            ch_rom[1318] <= 8'h00;
            ch_rom[1319] <= 8'h00;
            ch_rom[1320] <= 8'h00;
            ch_rom[1321] <= 8'h00;
            ch_rom[1322] <= 8'h00;
            ch_rom[1323] <= 8'h00;
            ch_rom[1324] <= 8'h00;
            ch_rom[1325] <= 8'h00;
            ch_rom[1326] <= 8'h00;
            ch_rom[1327] <= 8'h00;
            ch_rom[1328] <= 8'h00;
            ch_rom[1329] <= 8'h00;
            ch_rom[1330] <= 8'h00;
            ch_rom[1331] <= 8'h00;
            ch_rom[1332] <= 8'h00;
            ch_rom[1333] <= 8'h00;
            ch_rom[1334] <= 8'h00;
            ch_rom[1335] <= 8'h00;
            ch_rom[1336] <= 8'h00;
            ch_rom[1337] <= 8'h00;
            ch_rom[1338] <= 8'h00;
            ch_rom[1339] <= 8'h00;
            ch_rom[1340] <= 8'h00;
            ch_rom[1341] <= 8'h00;
            ch_rom[1342] <= 8'h00;
            ch_rom[1343] <= 8'h00;
            ch_rom[1344] <= 8'h00;
            ch_rom[1345] <= 8'h00;
            ch_rom[1346] <= 8'h00;
            ch_rom[1347] <= 8'h00;
            ch_rom[1348] <= 8'h00;
            ch_rom[1349] <= 8'h00;
            ch_rom[1350] <= 8'h00;
            ch_rom[1351] <= 8'h00;
            ch_rom[1352] <= 8'h00;
            ch_rom[1353] <= 8'h00;
            ch_rom[1354] <= 8'h00;
            ch_rom[1355] <= 8'h00;
            ch_rom[1356] <= 8'h00;
            ch_rom[1357] <= 8'h00;
            ch_rom[1358] <= 8'h00;
            ch_rom[1359] <= 8'h00;
            ch_rom[1360] <= 8'h00;
            ch_rom[1361] <= 8'h00;
            ch_rom[1362] <= 8'h00;
            ch_rom[1363] <= 8'h00;
            ch_rom[1364] <= 8'h00;
            ch_rom[1365] <= 8'h00;
            ch_rom[1366] <= 8'h00;
            ch_rom[1367] <= 8'h00;
            ch_rom[1368] <= 8'h00;
            ch_rom[1369] <= 8'h00;
            ch_rom[1370] <= 8'h00;
            ch_rom[1371] <= 8'h00;
            ch_rom[1372] <= 8'h00;
            ch_rom[1373] <= 8'h00;
            ch_rom[1374] <= 8'h00;
            ch_rom[1375] <= 8'h00;
            ch_rom[1376] <= 8'h00;
            ch_rom[1377] <= 8'h00;
            ch_rom[1378] <= 8'h00;
            ch_rom[1379] <= 8'h00;
            ch_rom[1380] <= 8'h00;
            ch_rom[1381] <= 8'h00;
            ch_rom[1382] <= 8'h00;
            ch_rom[1383] <= 8'h00;
            ch_rom[1384] <= 8'h00;
            ch_rom[1385] <= 8'h00;
            ch_rom[1386] <= 8'h00;
            ch_rom[1387] <= 8'h00;
            ch_rom[1388] <= 8'h00;
            ch_rom[1389] <= 8'h00;
            ch_rom[1390] <= 8'h00;
            ch_rom[1391] <= 8'h00;
            ch_rom[1392] <= 8'h00;
            ch_rom[1393] <= 8'h00;
            ch_rom[1394] <= 8'h00;
            ch_rom[1395] <= 8'h00;
            ch_rom[1396] <= 8'h00;
            ch_rom[1397] <= 8'h00;
            ch_rom[1398] <= 8'h00;
            ch_rom[1399] <= 8'h00;
            ch_rom[1400] <= 8'h00;
            ch_rom[1401] <= 8'h00;
            ch_rom[1402] <= 8'h00;
            ch_rom[1403] <= 8'h00;
            ch_rom[1404] <= 8'h00;
            ch_rom[1405] <= 8'h00;
            ch_rom[1406] <= 8'h00;
            ch_rom[1407] <= 8'h00;
            ch_rom[1408] <= 8'h00;
            ch_rom[1409] <= 8'h00;
            ch_rom[1410] <= 8'h00;
            ch_rom[1411] <= 8'h00;
            ch_rom[1412] <= 8'h00;
            ch_rom[1413] <= 8'h00;
            ch_rom[1414] <= 8'h00;
            ch_rom[1415] <= 8'h00;
            ch_rom[1416] <= 8'h00;
            ch_rom[1417] <= 8'h00;
            ch_rom[1418] <= 8'h00;
            ch_rom[1419] <= 8'h00;
            ch_rom[1420] <= 8'h00;
            ch_rom[1421] <= 8'h00;
            ch_rom[1422] <= 8'h00;
            ch_rom[1423] <= 8'h00;
            ch_rom[1424] <= 8'h00;
            ch_rom[1425] <= 8'h00;
            ch_rom[1426] <= 8'h00;
            ch_rom[1427] <= 8'h00;
            ch_rom[1428] <= 8'h00;
            ch_rom[1429] <= 8'h00;
            ch_rom[1430] <= 8'h00;
            ch_rom[1431] <= 8'h00;
            ch_rom[1432] <= 8'h00;
            ch_rom[1433] <= 8'h00;
            ch_rom[1434] <= 8'h00;
            ch_rom[1435] <= 8'h00;
            ch_rom[1436] <= 8'h00;
            ch_rom[1437] <= 8'h00;
            ch_rom[1438] <= 8'h00;
            ch_rom[1439] <= 8'h00;
            ch_rom[1440] <= 8'h00;
            ch_rom[1441] <= 8'h00;
            ch_rom[1442] <= 8'h00;
            ch_rom[1443] <= 8'h00;
            ch_rom[1444] <= 8'h00;
            ch_rom[1445] <= 8'h00;
            ch_rom[1446] <= 8'h00;
            ch_rom[1447] <= 8'h00;
            ch_rom[1448] <= 8'h00;
            ch_rom[1449] <= 8'h00;
            ch_rom[1450] <= 8'h00;
            ch_rom[1451] <= 8'h00;
            ch_rom[1452] <= 8'h00;
            ch_rom[1453] <= 8'h00;
            ch_rom[1454] <= 8'h00;
            ch_rom[1455] <= 8'h00;
            ch_rom[1456] <= 8'h00;
            ch_rom[1457] <= 8'h00;
            ch_rom[1458] <= 8'h00;
            ch_rom[1459] <= 8'h00;
            ch_rom[1460] <= 8'h00;
            ch_rom[1461] <= 8'h00;
            ch_rom[1462] <= 8'h00;
            ch_rom[1463] <= 8'h00;
            ch_rom[1464] <= 8'h00;
            ch_rom[1465] <= 8'h00;
            ch_rom[1466] <= 8'h00;
            ch_rom[1467] <= 8'h00;
            ch_rom[1468] <= 8'h00;
            ch_rom[1469] <= 8'h00;
            ch_rom[1470] <= 8'h00;
            ch_rom[1471] <= 8'h00;
            ch_rom[1472] <= 8'h00;
            ch_rom[1473] <= 8'h00;
            ch_rom[1474] <= 8'h00;
            ch_rom[1475] <= 8'h00;
            ch_rom[1476] <= 8'h00;
            ch_rom[1477] <= 8'h00;
            ch_rom[1478] <= 8'h00;
            ch_rom[1479] <= 8'h00;
            ch_rom[1480] <= 8'h00;
            ch_rom[1481] <= 8'h00;
            ch_rom[1482] <= 8'h00;
            ch_rom[1483] <= 8'h00;
            ch_rom[1484] <= 8'h00;
            ch_rom[1485] <= 8'h00;
            ch_rom[1486] <= 8'h00;
            ch_rom[1487] <= 8'h00;
            ch_rom[1488] <= 8'h00;
            ch_rom[1489] <= 8'h00;
            ch_rom[1490] <= 8'h00;
            ch_rom[1491] <= 8'h00;
            ch_rom[1492] <= 8'h00;
            ch_rom[1493] <= 8'h00;
            ch_rom[1494] <= 8'h00;
            ch_rom[1495] <= 8'h00;
            ch_rom[1496] <= 8'h00;
            ch_rom[1497] <= 8'h00;
            ch_rom[1498] <= 8'h00;
            ch_rom[1499] <= 8'h00;
            ch_rom[1500] <= 8'h00;
            ch_rom[1501] <= 8'h00;
            ch_rom[1502] <= 8'h00;
            ch_rom[1503] <= 8'h00;
            ch_rom[1504] <= 8'h00;
            ch_rom[1505] <= 8'h00;
            ch_rom[1506] <= 8'h00;
            ch_rom[1507] <= 8'h00;
            ch_rom[1508] <= 8'h00;
            ch_rom[1509] <= 8'h00;
            ch_rom[1510] <= 8'h00;
            ch_rom[1511] <= 8'h00;
            ch_rom[1512] <= 8'h00;
            ch_rom[1513] <= 8'h00;
            ch_rom[1514] <= 8'h00;
            ch_rom[1515] <= 8'h00;
            ch_rom[1516] <= 8'h00;
            ch_rom[1517] <= 8'h00;
            ch_rom[1518] <= 8'h00;
            ch_rom[1519] <= 8'h00;
            ch_rom[1520] <= 8'h00;
            ch_rom[1521] <= 8'h00;
            ch_rom[1522] <= 8'h00;
            ch_rom[1523] <= 8'h00;
            ch_rom[1524] <= 8'h00;
            ch_rom[1525] <= 8'h00;
            ch_rom[1526] <= 8'h00;
            ch_rom[1527] <= 8'h00;
            ch_rom[1528] <= 8'h00;
            ch_rom[1529] <= 8'h00;
            ch_rom[1530] <= 8'h00;
            ch_rom[1531] <= 8'h00;
            ch_rom[1532] <= 8'h00;
            ch_rom[1533] <= 8'h00;
            ch_rom[1534] <= 8'h00;
            ch_rom[1535] <= 8'h00;
            ch_rom[1536] <= 8'h00;
            ch_rom[1537] <= 8'h00;
            ch_rom[1538] <= 8'h00;
            ch_rom[1539] <= 8'h00;
            ch_rom[1540] <= 8'h00;
            ch_rom[1541] <= 8'h00;
            ch_rom[1542] <= 8'h00;
            ch_rom[1543] <= 8'h00;
            ch_rom[1544] <= 8'h00;
            ch_rom[1545] <= 8'h00;
            ch_rom[1546] <= 8'h00;
            ch_rom[1547] <= 8'h00;
            ch_rom[1548] <= 8'h00;
            ch_rom[1549] <= 8'h00;
            ch_rom[1550] <= 8'h00;
            ch_rom[1551] <= 8'h00;
            ch_rom[1552] <= 8'h00;
            ch_rom[1553] <= 8'h00;
            ch_rom[1554] <= 8'h00;
            ch_rom[1555] <= 8'h00;
            ch_rom[1556] <= 8'h00;
            ch_rom[1557] <= 8'h00;
            ch_rom[1558] <= 8'h00;
            ch_rom[1559] <= 8'h00;
            ch_rom[1560] <= 8'h00;
            ch_rom[1561] <= 8'h00;
            ch_rom[1562] <= 8'h00;
            ch_rom[1563] <= 8'h00;
            ch_rom[1564] <= 8'h00;
            ch_rom[1565] <= 8'h00;
            ch_rom[1566] <= 8'h00;
            ch_rom[1567] <= 8'h00;
            ch_rom[1568] <= 8'h00;
            ch_rom[1569] <= 8'h00;
            ch_rom[1570] <= 8'h00;
            ch_rom[1571] <= 8'h00;
            ch_rom[1572] <= 8'h00;
            ch_rom[1573] <= 8'h00;
            ch_rom[1574] <= 8'h00;
            ch_rom[1575] <= 8'h00;
            ch_rom[1576] <= 8'h00;
            ch_rom[1577] <= 8'h00;
            ch_rom[1578] <= 8'h00;
            ch_rom[1579] <= 8'h00;
            ch_rom[1580] <= 8'h00;
            ch_rom[1581] <= 8'h00;
            ch_rom[1582] <= 8'h00;
            ch_rom[1583] <= 8'h00;
            ch_rom[1584] <= 8'h00;
            ch_rom[1585] <= 8'h00;
            ch_rom[1586] <= 8'h00;
            ch_rom[1587] <= 8'h00;
            ch_rom[1588] <= 8'h00;
            ch_rom[1589] <= 8'h00;
            ch_rom[1590] <= 8'h00;
            ch_rom[1591] <= 8'h00;
            ch_rom[1592] <= 8'h00;
            ch_rom[1593] <= 8'h00;
            ch_rom[1594] <= 8'h00;
            ch_rom[1595] <= 8'h00;
            ch_rom[1596] <= 8'h00;
            ch_rom[1597] <= 8'h00;
            ch_rom[1598] <= 8'h00;
            ch_rom[1599] <= 8'h00;
            ch_rom[1600] <= 8'h00;
            ch_rom[1601] <= 8'h00;
            ch_rom[1602] <= 8'h00;
            ch_rom[1603] <= 8'h00;
            ch_rom[1604] <= 8'h00;
            ch_rom[1605] <= 8'h00;
            ch_rom[1606] <= 8'h00;
            ch_rom[1607] <= 8'h00;
            ch_rom[1608] <= 8'h00;
            ch_rom[1609] <= 8'h00;
            ch_rom[1610] <= 8'h00;
            ch_rom[1611] <= 8'h00;
            ch_rom[1612] <= 8'h00;
            ch_rom[1613] <= 8'h00;
            ch_rom[1614] <= 8'h00;
            ch_rom[1615] <= 8'h00;
            ch_rom[1616] <= 8'h00;
            ch_rom[1617] <= 8'h00;
            ch_rom[1618] <= 8'h00;
            ch_rom[1619] <= 8'h00;
            ch_rom[1620] <= 8'h00;
            ch_rom[1621] <= 8'h00;
            ch_rom[1622] <= 8'h00;
            ch_rom[1623] <= 8'h00;
            ch_rom[1624] <= 8'h00;
            ch_rom[1625] <= 8'h00;
            ch_rom[1626] <= 8'h00;
            ch_rom[1627] <= 8'h00;
            ch_rom[1628] <= 8'h00;
            ch_rom[1629] <= 8'h00;
            ch_rom[1630] <= 8'h00;
            ch_rom[1631] <= 8'h00;
            ch_rom[1632] <= 8'h00;
            ch_rom[1633] <= 8'h00;
            ch_rom[1634] <= 8'h00;
            ch_rom[1635] <= 8'h00;
            ch_rom[1636] <= 8'h00;
            ch_rom[1637] <= 8'h00;
            ch_rom[1638] <= 8'h00;
            ch_rom[1639] <= 8'h00;
            ch_rom[1640] <= 8'h00;
            ch_rom[1641] <= 8'h00;
            ch_rom[1642] <= 8'h00;
            ch_rom[1643] <= 8'h00;
            ch_rom[1644] <= 8'h00;
            ch_rom[1645] <= 8'h00;
            ch_rom[1646] <= 8'h00;
            ch_rom[1647] <= 8'h00;
            ch_rom[1648] <= 8'h00;
            ch_rom[1649] <= 8'h00;
            ch_rom[1650] <= 8'h00;
            ch_rom[1651] <= 8'h00;
            ch_rom[1652] <= 8'h00;
            ch_rom[1653] <= 8'h00;
            ch_rom[1654] <= 8'h00;
            ch_rom[1655] <= 8'h00;
            ch_rom[1656] <= 8'h00;
            ch_rom[1657] <= 8'h00;
            ch_rom[1658] <= 8'h00;
            ch_rom[1659] <= 8'h00;
            ch_rom[1660] <= 8'h00;
            ch_rom[1661] <= 8'h00;
            ch_rom[1662] <= 8'h00;
            ch_rom[1663] <= 8'h00;
            ch_rom[1664] <= 8'h00;
            ch_rom[1665] <= 8'h00;
            ch_rom[1666] <= 8'h00;
            ch_rom[1667] <= 8'h00;
            ch_rom[1668] <= 8'h00;
            ch_rom[1669] <= 8'h00;
            ch_rom[1670] <= 8'h00;
            ch_rom[1671] <= 8'h00;
            ch_rom[1672] <= 8'h00;
            ch_rom[1673] <= 8'h00;
            ch_rom[1674] <= 8'h00;
            ch_rom[1675] <= 8'h00;
            ch_rom[1676] <= 8'h00;
            ch_rom[1677] <= 8'h00;
            ch_rom[1678] <= 8'h00;
            ch_rom[1679] <= 8'h00;
            ch_rom[1680] <= 8'h00;
            ch_rom[1681] <= 8'h00;
            ch_rom[1682] <= 8'h00;
            ch_rom[1683] <= 8'h00;
            ch_rom[1684] <= 8'h00;
            ch_rom[1685] <= 8'h00;
            ch_rom[1686] <= 8'h00;
            ch_rom[1687] <= 8'h00;
            ch_rom[1688] <= 8'h00;
            ch_rom[1689] <= 8'h00;
            ch_rom[1690] <= 8'h00;
            ch_rom[1691] <= 8'h00;
            ch_rom[1692] <= 8'h00;
            ch_rom[1693] <= 8'h00;
            ch_rom[1694] <= 8'h00;
            ch_rom[1695] <= 8'h00;
            ch_rom[1696] <= 8'h00;
            ch_rom[1697] <= 8'h00;
            ch_rom[1698] <= 8'h00;
            ch_rom[1699] <= 8'h00;
            ch_rom[1700] <= 8'h00;
            ch_rom[1701] <= 8'h00;
            ch_rom[1702] <= 8'h00;
            ch_rom[1703] <= 8'h00;
            ch_rom[1704] <= 8'h00;
            ch_rom[1705] <= 8'h00;
            ch_rom[1706] <= 8'h00;
            ch_rom[1707] <= 8'h00;
            ch_rom[1708] <= 8'h00;
            ch_rom[1709] <= 8'h00;
            ch_rom[1710] <= 8'h00;
            ch_rom[1711] <= 8'h00;
            ch_rom[1712] <= 8'h00;
            ch_rom[1713] <= 8'h00;
            ch_rom[1714] <= 8'h00;
            ch_rom[1715] <= 8'h00;
            ch_rom[1716] <= 8'h00;
            ch_rom[1717] <= 8'h00;
            ch_rom[1718] <= 8'h00;
            ch_rom[1719] <= 8'h00;
            ch_rom[1720] <= 8'h00;
            ch_rom[1721] <= 8'h00;
            ch_rom[1722] <= 8'h00;
            ch_rom[1723] <= 8'h00;
            ch_rom[1724] <= 8'h00;
            ch_rom[1725] <= 8'h00;
            ch_rom[1726] <= 8'h00;
            ch_rom[1727] <= 8'h00;
            ch_rom[1728] <= 8'h00;
            ch_rom[1729] <= 8'h00;
            ch_rom[1730] <= 8'h00;
            ch_rom[1731] <= 8'h00;
            ch_rom[1732] <= 8'h00;
            ch_rom[1733] <= 8'h00;
            ch_rom[1734] <= 8'h00;
            ch_rom[1735] <= 8'h00;
            ch_rom[1736] <= 8'h00;
            ch_rom[1737] <= 8'h00;
            ch_rom[1738] <= 8'h00;
            ch_rom[1739] <= 8'h00;
            ch_rom[1740] <= 8'h00;
            ch_rom[1741] <= 8'h00;
            ch_rom[1742] <= 8'h00;
            ch_rom[1743] <= 8'h00;
            ch_rom[1744] <= 8'h00;
            ch_rom[1745] <= 8'h00;
            ch_rom[1746] <= 8'h00;
            ch_rom[1747] <= 8'h00;
            ch_rom[1748] <= 8'h00;
            ch_rom[1749] <= 8'h00;
            ch_rom[1750] <= 8'h00;
            ch_rom[1751] <= 8'h00;
            ch_rom[1752] <= 8'h00;
            ch_rom[1753] <= 8'h00;
            ch_rom[1754] <= 8'h00;
            ch_rom[1755] <= 8'h00;
            ch_rom[1756] <= 8'h00;
            ch_rom[1757] <= 8'h00;
            ch_rom[1758] <= 8'h00;
            ch_rom[1759] <= 8'h00;
            ch_rom[1760] <= 8'h00;
            ch_rom[1761] <= 8'h00;
            ch_rom[1762] <= 8'h00;
            ch_rom[1763] <= 8'h00;
            ch_rom[1764] <= 8'h00;
            ch_rom[1765] <= 8'h00;
            ch_rom[1766] <= 8'h00;
            ch_rom[1767] <= 8'h00;
            ch_rom[1768] <= 8'h00;
            ch_rom[1769] <= 8'h00;
            ch_rom[1770] <= 8'h00;
            ch_rom[1771] <= 8'h00;
            ch_rom[1772] <= 8'h00;
            ch_rom[1773] <= 8'h00;
            ch_rom[1774] <= 8'h00;
            ch_rom[1775] <= 8'h00;
            ch_rom[1776] <= 8'h00;
            ch_rom[1777] <= 8'h00;
            ch_rom[1778] <= 8'h00;
            ch_rom[1779] <= 8'h00;
            ch_rom[1780] <= 8'h00;
            ch_rom[1781] <= 8'h00;
            ch_rom[1782] <= 8'h00;
            ch_rom[1783] <= 8'h00;
            ch_rom[1784] <= 8'h00;
            ch_rom[1785] <= 8'h00;
            ch_rom[1786] <= 8'h00;
            ch_rom[1787] <= 8'h00;
            ch_rom[1788] <= 8'h00;
            ch_rom[1789] <= 8'h00;
            ch_rom[1790] <= 8'h00;
            ch_rom[1791] <= 8'h00;
            ch_rom[1792] <= 8'h00;
            ch_rom[1793] <= 8'h00;
            ch_rom[1794] <= 8'h00;
            ch_rom[1795] <= 8'h00;
            ch_rom[1796] <= 8'h00;
            ch_rom[1797] <= 8'h00;
            ch_rom[1798] <= 8'h00;
            ch_rom[1799] <= 8'h00;
            ch_rom[1800] <= 8'h00;
            ch_rom[1801] <= 8'h00;
            ch_rom[1802] <= 8'h00;
            ch_rom[1803] <= 8'h00;
            ch_rom[1804] <= 8'h00;
            ch_rom[1805] <= 8'h00;
            ch_rom[1806] <= 8'h00;
            ch_rom[1807] <= 8'h00;
            ch_rom[1808] <= 8'h00;
            ch_rom[1809] <= 8'h00;
            ch_rom[1810] <= 8'h00;
            ch_rom[1811] <= 8'h00;
            ch_rom[1812] <= 8'h00;
            ch_rom[1813] <= 8'h00;
            ch_rom[1814] <= 8'h00;
            ch_rom[1815] <= 8'h00;
            ch_rom[1816] <= 8'h00;
            ch_rom[1817] <= 8'h00;
            ch_rom[1818] <= 8'h00;
            ch_rom[1819] <= 8'h00;
            ch_rom[1820] <= 8'h00;
            ch_rom[1821] <= 8'h00;
            ch_rom[1822] <= 8'h00;
            ch_rom[1823] <= 8'h00;
            ch_rom[1824] <= 8'h00;
            ch_rom[1825] <= 8'h00;
            ch_rom[1826] <= 8'h00;
            ch_rom[1827] <= 8'h00;
            ch_rom[1828] <= 8'h00;
            ch_rom[1829] <= 8'h00;
            ch_rom[1830] <= 8'h00;
            ch_rom[1831] <= 8'h00;
            ch_rom[1832] <= 8'h00;
            ch_rom[1833] <= 8'h00;
            ch_rom[1834] <= 8'h00;
            ch_rom[1835] <= 8'h00;
            ch_rom[1836] <= 8'h00;
            ch_rom[1837] <= 8'h00;
            ch_rom[1838] <= 8'h00;
            ch_rom[1839] <= 8'h00;
            ch_rom[1840] <= 8'h00;
            ch_rom[1841] <= 8'h00;
            ch_rom[1842] <= 8'h00;
            ch_rom[1843] <= 8'h00;
            ch_rom[1844] <= 8'h00;
            ch_rom[1845] <= 8'h00;
            ch_rom[1846] <= 8'h00;
            ch_rom[1847] <= 8'h00;
            ch_rom[1848] <= 8'h00;
            ch_rom[1849] <= 8'h00;
            ch_rom[1850] <= 8'h00;
            ch_rom[1851] <= 8'h00;
            ch_rom[1852] <= 8'h00;
            ch_rom[1853] <= 8'h00;
            ch_rom[1854] <= 8'h00;
            ch_rom[1855] <= 8'h00;
            ch_rom[1856] <= 8'h00;
            ch_rom[1857] <= 8'h00;
            ch_rom[1858] <= 8'h00;
            ch_rom[1859] <= 8'h00;
            ch_rom[1860] <= 8'h00;
            ch_rom[1861] <= 8'h00;
            ch_rom[1862] <= 8'h00;
            ch_rom[1863] <= 8'h00;
            ch_rom[1864] <= 8'h00;
            ch_rom[1865] <= 8'h00;
            ch_rom[1866] <= 8'h00;
            ch_rom[1867] <= 8'h00;
            ch_rom[1868] <= 8'h00;
            ch_rom[1869] <= 8'h00;
            ch_rom[1870] <= 8'h00;
            ch_rom[1871] <= 8'h00;
            ch_rom[1872] <= 8'h00;
            ch_rom[1873] <= 8'h00;
            ch_rom[1874] <= 8'h00;
            ch_rom[1875] <= 8'h00;
            ch_rom[1876] <= 8'h00;
            ch_rom[1877] <= 8'h00;
            ch_rom[1878] <= 8'h00;
            ch_rom[1879] <= 8'h00;
            ch_rom[1880] <= 8'h00;
            ch_rom[1881] <= 8'h00;
            ch_rom[1882] <= 8'h00;
            ch_rom[1883] <= 8'h00;
            ch_rom[1884] <= 8'h00;
            ch_rom[1885] <= 8'h00;
            ch_rom[1886] <= 8'h00;
            ch_rom[1887] <= 8'h00;
            ch_rom[1888] <= 8'h00;
            ch_rom[1889] <= 8'h00;
            ch_rom[1890] <= 8'h00;
            ch_rom[1891] <= 8'h00;
            ch_rom[1892] <= 8'h00;
            ch_rom[1893] <= 8'h00;
            ch_rom[1894] <= 8'h00;
            ch_rom[1895] <= 8'h00;
            ch_rom[1896] <= 8'h00;
            ch_rom[1897] <= 8'h00;
            ch_rom[1898] <= 8'h00;
            ch_rom[1899] <= 8'h00;
            ch_rom[1900] <= 8'h00;
            ch_rom[1901] <= 8'h00;
            ch_rom[1902] <= 8'h00;
            ch_rom[1903] <= 8'h00;
            ch_rom[1904] <= 8'h00;
            ch_rom[1905] <= 8'h00;
            ch_rom[1906] <= 8'h00;
            ch_rom[1907] <= 8'h00;
            ch_rom[1908] <= 8'h00;
            ch_rom[1909] <= 8'h00;
            ch_rom[1910] <= 8'h00;
            ch_rom[1911] <= 8'h00;
            ch_rom[1912] <= 8'h00;
            ch_rom[1913] <= 8'h00;
            ch_rom[1914] <= 8'h00;
            ch_rom[1915] <= 8'h00;
            ch_rom[1916] <= 8'h00;
            ch_rom[1917] <= 8'h00;
            ch_rom[1918] <= 8'h00;
            ch_rom[1919] <= 8'h00;
            ch_rom[1920] <= 8'h00;
            ch_rom[1921] <= 8'h00;
            ch_rom[1922] <= 8'h00;
            ch_rom[1923] <= 8'h00;
            ch_rom[1924] <= 8'h00;
            ch_rom[1925] <= 8'h00;
            ch_rom[1926] <= 8'h00;
            ch_rom[1927] <= 8'h00;
            ch_rom[1928] <= 8'h00;
            ch_rom[1929] <= 8'h00;
            ch_rom[1930] <= 8'h00;
            ch_rom[1931] <= 8'h00;
            ch_rom[1932] <= 8'h00;
            ch_rom[1933] <= 8'h00;
            ch_rom[1934] <= 8'h00;
            ch_rom[1935] <= 8'h00;
            ch_rom[1936] <= 8'h00;
            ch_rom[1937] <= 8'h00;
            ch_rom[1938] <= 8'h00;
            ch_rom[1939] <= 8'h00;
            ch_rom[1940] <= 8'h00;
            ch_rom[1941] <= 8'h00;
            ch_rom[1942] <= 8'h00;
            ch_rom[1943] <= 8'h00;
            ch_rom[1944] <= 8'h00;
            ch_rom[1945] <= 8'h00;
            ch_rom[1946] <= 8'h00;
            ch_rom[1947] <= 8'h00;
            ch_rom[1948] <= 8'h00;
            ch_rom[1949] <= 8'h00;
            ch_rom[1950] <= 8'h00;
            ch_rom[1951] <= 8'h00;
            ch_rom[1952] <= 8'h00;
            ch_rom[1953] <= 8'h00;
            ch_rom[1954] <= 8'h00;
            ch_rom[1955] <= 8'h00;
            ch_rom[1956] <= 8'h00;
            ch_rom[1957] <= 8'h00;
            ch_rom[1958] <= 8'h00;
            ch_rom[1959] <= 8'h00;
            ch_rom[1960] <= 8'h00;
            ch_rom[1961] <= 8'h00;
            ch_rom[1962] <= 8'h00;
            ch_rom[1963] <= 8'h00;
            ch_rom[1964] <= 8'h00;
            ch_rom[1965] <= 8'h00;
            ch_rom[1966] <= 8'h00;
            ch_rom[1967] <= 8'h00;
            ch_rom[1968] <= 8'h00;
            ch_rom[1969] <= 8'h00;
            ch_rom[1970] <= 8'h00;
            ch_rom[1971] <= 8'h00;
            ch_rom[1972] <= 8'h00;
            ch_rom[1973] <= 8'h00;
            ch_rom[1974] <= 8'h00;
            ch_rom[1975] <= 8'h00;
            ch_rom[1976] <= 8'h00;
            ch_rom[1977] <= 8'h00;
            ch_rom[1978] <= 8'h00;
            ch_rom[1979] <= 8'h00;
            ch_rom[1980] <= 8'h00;
            ch_rom[1981] <= 8'h00;
            ch_rom[1982] <= 8'h00;
            ch_rom[1983] <= 8'h00;
            ch_rom[1984] <= 8'h00;
            ch_rom[1985] <= 8'h00;
            ch_rom[1986] <= 8'h00;
            ch_rom[1987] <= 8'h00;
            ch_rom[1988] <= 8'h00;
            ch_rom[1989] <= 8'h00;
            ch_rom[1990] <= 8'h00;
            ch_rom[1991] <= 8'h00;
            ch_rom[1992] <= 8'h00;
            ch_rom[1993] <= 8'h00;
            ch_rom[1994] <= 8'h00;
            ch_rom[1995] <= 8'h00;
            ch_rom[1996] <= 8'h00;
            ch_rom[1997] <= 8'h00;
            ch_rom[1998] <= 8'h00;
            ch_rom[1999] <= 8'h00;
            ch_rom[2000] <= 8'h00;
            ch_rom[2001] <= 8'h00;
            ch_rom[2002] <= 8'h00;
            ch_rom[2003] <= 8'h00;
            ch_rom[2004] <= 8'h00;
            ch_rom[2005] <= 8'h00;
            ch_rom[2006] <= 8'h00;
            ch_rom[2007] <= 8'h00;
            ch_rom[2008] <= 8'h00;
            ch_rom[2009] <= 8'h00;
            ch_rom[2010] <= 8'h00;
            ch_rom[2011] <= 8'h00;
            ch_rom[2012] <= 8'h00;
            ch_rom[2013] <= 8'h00;
            ch_rom[2014] <= 8'h00;
            ch_rom[2015] <= 8'h00;
            ch_rom[2016] <= 8'h00;
            ch_rom[2017] <= 8'h00;
            ch_rom[2018] <= 8'h00;
            ch_rom[2019] <= 8'h00;
            ch_rom[2020] <= 8'h00;
            ch_rom[2021] <= 8'h00;
            ch_rom[2022] <= 8'h00;
            ch_rom[2023] <= 8'h00;
            ch_rom[2024] <= 8'h00;
            ch_rom[2025] <= 8'h00;
            ch_rom[2026] <= 8'h00;
            ch_rom[2027] <= 8'h00;
            ch_rom[2028] <= 8'h00;
            ch_rom[2029] <= 8'h00;
            ch_rom[2030] <= 8'h00;
            ch_rom[2031] <= 8'h00;
            ch_rom[2032] <= 8'h00;
            ch_rom[2033] <= 8'h00;
            ch_rom[2034] <= 8'h00;
            ch_rom[2035] <= 8'h00;
            ch_rom[2036] <= 8'h00;
            ch_rom[2037] <= 8'h00;
            ch_rom[2038] <= 8'h00;
            ch_rom[2039] <= 8'h00;
            ch_rom[2040] <= 8'h00;
            ch_rom[2041] <= 8'h00;
            ch_rom[2042] <= 8'h00;
            ch_rom[2043] <= 8'h00;
            ch_rom[2044] <= 8'h00;
            ch_rom[2045] <= 8'h00;
            ch_rom[2046] <= 8'h00;
            ch_rom[2047] <= 8'h00;
        end
    end
endmodule
